// Given a board state, return the move that X should make.
`default_nettype none
module xmove(i_board, o_move);
  input wire [17:0] i_board;
  output reg [3:0]  o_move;

  always @(*) 
    case (i_board)
      18'b010001011100110000: begin o_move = 4'd2; end
      18'b010100011100110000: begin o_move = 4'd3; end
      18'b000001011101000011: begin o_move = 4'd1; end
      18'b000101001101000011: begin o_move = 4'd1; end
      18'b010000011101110000: begin o_move = 4'd2; end
      18'b010001001101000011: begin o_move = 4'd2; end
      18'b010111011100000000: begin o_move = 4'd7; end
      18'b000001011100000000: begin o_move = 4'd1; end
      18'b000101001100000000: begin o_move = 4'd1; end
      18'b010001001100000000: begin o_move = 4'd2; end
      18'b010100001100000000: begin o_move = 4'd3; end
      18'b010000011100000000: begin o_move = 4'd7; end
      18'b000101111101000111: begin o_move = 4'd1; end
      18'b010001111101000111: begin o_move = 4'd2; end
      18'b010001111100010111: begin o_move = 4'd6; end
      18'b010100111100010111: begin o_move = 4'd6; end
      18'b010111110101000011: begin o_move = 4'd8; end
      18'b010111110101001100: begin o_move = 4'd9; end
      18'b000001011111000001: begin o_move = 4'd1; end
      18'b000101111100000100: begin o_move = 4'd1; end
      18'b010000011100110001: begin o_move = 4'd2; end
      18'b010001001111000001: begin o_move = 4'd2; end
      18'b010001111100010000: begin o_move = 4'd2; end
      18'b010000011100110100: begin o_move = 4'd3; end
      18'b010100111100000100: begin o_move = 4'd3; end
      18'b000101001111000001: begin o_move = 4'd4; end
      18'b010111001100000001: begin o_move = 4'd4; end
      18'b010111001100000100: begin o_move = 4'd4; end
      18'b010111001100010000: begin o_move = 4'd4; end
      18'b010111110001000000: begin o_move = 4'd5; end
      18'b010001111100000100: begin o_move = 4'd6; end
      18'b010100111100010000: begin o_move = 4'd6; end
      18'b010111001101000000: begin o_move = 4'd7; end
      18'b010111110001110001: begin o_move = 4'd5; end
      18'b000001011111110101: begin o_move = 4'd1; end
      18'b000101001111110101: begin o_move = 4'd4; end
      18'b010001001111110101: begin o_move = 4'd4; end
      18'b010111111100000101: begin o_move = 4'd6; end
      18'b010111111100010001: begin o_move = 4'd6; end
      18'b010111111100010100: begin o_move = 4'd6; end
      18'b010111111101000001: begin o_move = 4'd7; end
      18'b010111111101000100: begin o_move = 4'd7; end
      18'b010111111101010000: begin o_move = 4'd8; end
      18'b000000000100000000: begin o_move = 4'd1; end
      18'b000000010000000000: begin o_move = 4'd1; end
      18'b000100000000000000: begin o_move = 4'd1; end
      18'b000000000000000100: begin o_move = 4'd2; end
      18'b000000000001000000: begin o_move = 4'd3; end
      18'b000000000000000001: begin o_move = 4'd5; end
      18'b000000000000010000: begin o_move = 4'd5; end
      18'b000001000000000000: begin o_move = 4'd5; end
      18'b010000000000000000: begin o_move = 4'd5; end
      18'b011100000101110111: begin o_move = 4'd4; end
      18'b011101000001110111: begin o_move = 4'd4; end
      18'b011101000100110111: begin o_move = 4'd4; end
      18'b011100010100110111: begin o_move = 4'd6; end
      18'b011101011101000011: begin o_move = 4'd8; end
      18'b011101011101110000: begin o_move = 4'd8; end
      18'b000000011100010111: begin o_move = 4'd1; end
      18'b000001001100010111: begin o_move = 4'd1; end
      18'b000001001101000111: begin o_move = 4'd1; end
      18'b000001001101010011: begin o_move = 4'd1; end
      18'b000100001100010111: begin o_move = 4'd1; end
      18'b010000001100010111: begin o_move = 4'd4; end
      18'b011100000000010111: begin o_move = 4'd4; end
      18'b011101011100000000: begin o_move = 4'd8; end
      18'b011101011100110100: begin o_move = 4'd6; end
      18'b011101011100110001: begin o_move = 4'd8; end
      18'b011101011111000001: begin o_move = 4'd8; end
      18'b011100010111110100: begin o_move = 4'd9; end
      18'b000000011100000001: begin o_move = 4'd1; end
      18'b000000011100010000: begin o_move = 4'd1; end
      18'b000100001100000001: begin o_move = 4'd1; end
      18'b000100001100010000: begin o_move = 4'd1; end
      18'b000001001100010000: begin o_move = 4'd2; end
      18'b010000001100000001: begin o_move = 4'd2; end
      18'b010000001101000000: begin o_move = 4'd2; end
      18'b000001001100000100: begin o_move = 4'd4; end
      18'b000111000001000000: begin o_move = 4'd4; end
      18'b010000001100000100: begin o_move = 4'd4; end
      18'b010000001100010000: begin o_move = 4'd4; end
      18'b010011000001000000: begin o_move = 4'd4; end
      18'b000001001100000001: begin o_move = 4'd6; end
      18'b011100000000000100: begin o_move = 4'd7; end
      18'b000001001101000000: begin o_move = 4'd9; end
      18'b011101001100010111: begin o_move = 4'd4; end
      18'b011101001101000111: begin o_move = 4'd4; end
      18'b011101110000010111: begin o_move = 4'd5; end
      18'b011101001101010011: begin o_move = 4'd8; end
      18'b000100001100011101: begin o_move = 4'd1; end
      18'b000111011101000000: begin o_move = 4'd1; end
      18'b000000011100011101: begin o_move = 4'd2; end
      18'b000001001100011101: begin o_move = 4'd2; end
      18'b010000001100011101: begin o_move = 4'd2; end
      18'b011101001100000100: begin o_move = 4'd4; end
      18'b011101001100010000: begin o_move = 4'd4; end
      18'b011100000001110100: begin o_move = 4'd5; end
      18'b011100010000110100: begin o_move = 4'd5; end
      18'b011101000000110100: begin o_move = 4'd5; end
      18'b011101001100000001: begin o_move = 4'd6; end
      18'b010011011101000000: begin o_move = 4'd7; end
      18'b011100011100000001: begin o_move = 4'd7; end
      18'b011100011101000000: begin o_move = 4'd7; end
      18'b011101001101000000: begin o_move = 4'd8; end
      18'b011100000100110100: begin o_move = 4'd9; end
      18'b011100011101110001: begin o_move = 4'd3; end
      18'b011100011101110100: begin o_move = 4'd3; end
      18'b011101001101110100: begin o_move = 4'd9; end
      18'b011100011100110101: begin o_move = 4'd3; end
      18'b011101001111000101: begin o_move = 4'd4; end
      18'b011101001111010001: begin o_move = 4'd4; end
      18'b011101000011110101: begin o_move = 4'd5; end
      18'b011101001100110101: begin o_move = 4'd6; end
      18'b011101111100000101: begin o_move = 4'd6; end
      18'b011101111100010001: begin o_move = 4'd6; end
      18'b011101111100010100: begin o_move = 4'd6; end
      18'b011101111101010000: begin o_move = 4'd8; end
      18'b011101111101000100: begin o_move = 4'd9; end
      18'b000001111101010111: begin o_move = 4'd1; end
      18'b000111110101011100: begin o_move = 4'd1; end
      18'b010000111101010111: begin o_move = 4'd2; end
      18'b010011110101000111: begin o_move = 4'd2; end
      18'b010011110101010011: begin o_move = 4'd2; end
      18'b011100110001010111: begin o_move = 4'd3; end
      18'b011100110100010111: begin o_move = 4'd3; end
      18'b011100001101010111: begin o_move = 4'd4; end
      18'b011111000100010111: begin o_move = 4'd6; end
      18'b000100001100110101: begin o_move = 4'd1; end
      18'b010000111101010000: begin o_move = 4'd2; end
      18'b010011001101000001: begin o_move = 4'd2; end
      18'b000000011100110101: begin o_move = 4'd3; end
      18'b010000001100110101: begin o_move = 4'd3; end
      18'b010000111101000100: begin o_move = 4'd3; end
      18'b011100001101000001: begin o_move = 4'd3; end
      18'b000001001111000101: begin o_move = 4'd4; end
      18'b000001001111010001: begin o_move = 4'd4; end
      18'b000111110001000100: begin o_move = 4'd5; end
      18'b000111110001010000: begin o_move = 4'd5; end
      18'b010011110001000001: begin o_move = 4'd5; end
      18'b010011110001000100: begin o_move = 4'd5; end
      18'b010011110001010000: begin o_move = 4'd5; end
      18'b011100000000110101: begin o_move = 4'd5; end
      18'b000001001100110101: begin o_move = 4'd6; end
      18'b000001111100000101: begin o_move = 4'd6; end
      18'b000001111100010100: begin o_move = 4'd6; end
      18'b010000111100000101: begin o_move = 4'd6; end
      18'b010000111100010001: begin o_move = 4'd6; end
      18'b010000111100010100: begin o_move = 4'd6; end
      18'b000111001101000001: begin o_move = 4'd7; end
      18'b000111110001000001: begin o_move = 4'd7; end
      18'b011100001100000101: begin o_move = 4'd7; end
      18'b011100001101000100: begin o_move = 4'd7; end
      18'b000111110101000000: begin o_move = 4'd8; end
      18'b011100001100010001: begin o_move = 4'd8; end
      18'b011100001101010000: begin o_move = 4'd8; end
      18'b000001111101000100: begin o_move = 4'd9; end
      18'b010011110101000000: begin o_move = 4'd9; end
      18'b000111001101011101: begin o_move = 4'd1; end
      18'b000111110101001101: begin o_move = 4'd1; end
      18'b000111110101110001: begin o_move = 4'd1; end
      18'b010011001101011101: begin o_move = 4'd2; end
      18'b011100110101110100: begin o_move = 4'd9; end
      18'b000111110001110101: begin o_move = 4'd1; end
      18'b011100001101110101: begin o_move = 4'd3; end
      18'b011111000001110101: begin o_move = 4'd5; end
      18'b011111010000110101: begin o_move = 4'd5; end
      18'b011111011101000001: begin o_move = 4'd7; end
      18'b000111111101000101: begin o_move = 4'd7; end
      18'b010011111101000101: begin o_move = 4'd7; end
      18'b011111001101000101: begin o_move = 4'd7; end
      18'b000111111101010001: begin o_move = 4'd8; end
      18'b010011111101010001: begin o_move = 4'd8; end
      18'b011100111101010001: begin o_move = 4'd8; end
      18'b011111001101010001: begin o_move = 4'd8; end
      18'b000111111101010100: begin o_move = 4'd9; end
      18'b010011111101010100: begin o_move = 4'd9; end
      18'b011100111101010100: begin o_move = 4'd9; end
      18'b011111110101000100: begin o_move = 4'd9; end
      18'b110101000101111100: begin o_move = 4'd4; end
      18'b110101010111001100: begin o_move = 4'd7; end
      18'b110101010111110000: begin o_move = 4'd8; end
      18'b110101010100111100: begin o_move = 4'd9; end
      18'b110100010111011100: begin o_move = 4'd3; end
      18'b001101000101110111: begin o_move = 4'd4; end
      18'b001101010001110111: begin o_move = 4'd5; end
      18'b110101011101110000: begin o_move = 4'd9; end
      18'b000000001101010111: begin o_move = 4'd1; end
      18'b001100000001010111: begin o_move = 4'd1; end
      18'b001100010000010111: begin o_move = 4'd1; end
      18'b001100000100010111: begin o_move = 4'd3; end
      18'b110100000100011100: begin o_move = 4'd3; end
      18'b110001000101110000: begin o_move = 4'd4; end
      18'b110100000101001100: begin o_move = 4'd4; end
      18'b110100000101110000: begin o_move = 4'd4; end
      18'b110101000001110000: begin o_move = 4'd4; end
      18'b110101000100110000: begin o_move = 4'd4; end
      18'b001101000000010111: begin o_move = 4'd5; end
      18'b110100010001110000: begin o_move = 4'd5; end
      18'b110001010100110000: begin o_move = 4'd6; end
      18'b110100010100001100: begin o_move = 4'd6; end
      18'b110001010111000000: begin o_move = 4'd7; end
      18'b110101000100001100: begin o_move = 4'd7; end
      18'b110100010111000000: begin o_move = 4'd8; end
      18'b110101011100000000: begin o_move = 4'd9; end
      18'b001101010111110100: begin o_move = 4'd1; end
      18'b110001010111110001: begin o_move = 4'd2; end
      18'b110001010111110100: begin o_move = 4'd2; end
      18'b110100010111001101: begin o_move = 4'd3; end
      18'b110101000100111101: begin o_move = 4'd4; end
      18'b110101011111000001: begin o_move = 4'd7; end
      18'b000011000001000001: begin o_move = 4'd1; end
      18'b000011000001000100: begin o_move = 4'd1; end
      18'b000011000001010000: begin o_move = 4'd1; end
      18'b001100000100000100: begin o_move = 4'd1; end
      18'b000000001101010000: begin o_move = 4'd2; end
      18'b110000000100000100: begin o_move = 4'd2; end
      18'b110000010000010000: begin o_move = 4'd2; end
      18'b000000001101000001: begin o_move = 4'd3; end
      18'b110000000100000001: begin o_move = 4'd3; end
      18'b110000000100010000: begin o_move = 4'd3; end
      18'b110000010000000001: begin o_move = 4'd3; end
      18'b110000010000000100: begin o_move = 4'd3; end
      18'b000011000101000000: begin o_move = 4'd4; end
      18'b110000000101000000: begin o_move = 4'd4; end
      18'b110101000000000000: begin o_move = 4'd4; end
      18'b000011010001000000: begin o_move = 4'd5; end
      18'b110000010001000000: begin o_move = 4'd5; end
      18'b110001010000000000: begin o_move = 4'd5; end
      18'b110100000000000001: begin o_move = 4'd5; end
      18'b110100000000000100: begin o_move = 4'd5; end
      18'b110100000000010000: begin o_move = 4'd5; end
      18'b110100010000000000: begin o_move = 4'd5; end
      18'b110000010100000000: begin o_move = 4'd6; end
      18'b000000001100000101: begin o_move = 4'd7; end
      18'b001100000000000101: begin o_move = 4'd7; end
      18'b001100000001000100: begin o_move = 4'd7; end
      18'b001100010000000100: begin o_move = 4'd7; end
      18'b001101000000000100: begin o_move = 4'd7; end
      18'b110001000100000000: begin o_move = 4'd7; end
      18'b110100000001000000: begin o_move = 4'd7; end
      18'b000000001100010001: begin o_move = 4'd8; end
      18'b110100000100000000: begin o_move = 4'd8; end
      18'b000000001100010100: begin o_move = 4'd9; end
      18'b001100000000010100: begin o_move = 4'd9; end
      18'b001101011100010111: begin o_move = 4'd1; end
      18'b110101110101001100: begin o_move = 4'd7; end
      18'b001101000100110100: begin o_move = 4'd1; end
      18'b001101011100010000: begin o_move = 4'd1; end
      18'b000000001101011101: begin o_move = 4'd2; end
      18'b110000010111000001: begin o_move = 4'd2; end
      18'b110000010111000100: begin o_move = 4'd2; end
      18'b110001011100010000: begin o_move = 4'd2; end
      18'b110000010111010000: begin o_move = 4'd3; end
      18'b110100000001110001: begin o_move = 4'd3; end
      18'b110100000100001101: begin o_move = 4'd3; end
      18'b110100011100000001: begin o_move = 4'd3; end
      18'b110100011100000100: begin o_move = 4'd3; end
      18'b110100011101000000: begin o_move = 4'd3; end
      18'b001100000101110100: begin o_move = 4'd4; end
      18'b110001000100110001: begin o_move = 4'd4; end
      18'b110001000100110100: begin o_move = 4'd4; end
      18'b110100000001110100: begin o_move = 4'd4; end
      18'b110101001100000100: begin o_move = 4'd4; end
      18'b110101001100010000: begin o_move = 4'd4; end
      18'b001100010001110100: begin o_move = 4'd5; end
      18'b001101010000110100: begin o_move = 4'd5; end
      18'b110101110000000100: begin o_move = 4'd5; end
      18'b110101110000010000: begin o_move = 4'd5; end
      18'b001100010100110100: begin o_move = 4'd6; end
      18'b110001011100000001: begin o_move = 4'd6; end
      18'b110101001100000001: begin o_move = 4'd6; end
      18'b110101110000000001: begin o_move = 4'd6; end
      18'b110101110001000000: begin o_move = 4'd7; end
      18'b110101110100000000: begin o_move = 4'd7; end
      18'b001101000001110100: begin o_move = 4'd9; end
      18'b110001011100000100: begin o_move = 4'd9; end
      18'b110001011101000000: begin o_move = 4'd9; end
      18'b110100011100010000: begin o_move = 4'd9; end
      18'b110101001101000000: begin o_move = 4'd9; end
      18'b110001011100011101: begin o_move = 4'd2; end
      18'b110100011100011101: begin o_move = 4'd3; end
      18'b110100011101110001: begin o_move = 4'd3; end
      18'b110100011101110100: begin o_move = 4'd3; end
      18'b110101001100011101: begin o_move = 4'd6; end
      18'b110101110111000001: begin o_move = 4'd7; end
      18'b001101011101110100: begin o_move = 4'd9; end
      18'b001100010111110101: begin o_move = 4'd1; end
      18'b001101000111110101: begin o_move = 4'd1; end
      18'b001101010011110101: begin o_move = 4'd1; end
      18'b110100011100110101: begin o_move = 4'd3; end
      18'b110101001100110101: begin o_move = 4'd4; end
      18'b110101001111000101: begin o_move = 4'd4; end
      18'b110101001111010001: begin o_move = 4'd4; end
      18'b110101110011000101: begin o_move = 4'd5; end
      18'b110101110011010001: begin o_move = 4'd5; end
      18'b001101011100110101: begin o_move = 4'd6; end
      18'b110001011100110101: begin o_move = 4'd6; end
      18'b110101111100000101: begin o_move = 4'd6; end
      18'b110101111100010001: begin o_move = 4'd6; end
      18'b110101111100010100: begin o_move = 4'd6; end
      18'b110001011111000101: begin o_move = 4'd7; end
      18'b110101111101000100: begin o_move = 4'd7; end
      18'b110001011111010001: begin o_move = 4'd8; end
      18'b110101111101010000: begin o_move = 4'd9; end
      18'b001100011101010111: begin o_move = 4'd1; end
      18'b001101001101010111: begin o_move = 4'd1; end
      18'b110100110101011100: begin o_move = 4'd3; end
      18'b110111000101011100: begin o_move = 4'd4; end
      18'b110111010100011100: begin o_move = 4'd6; end
      18'b000011011101000001: begin o_move = 4'd1; end
      18'b000011011101000100: begin o_move = 4'd1; end
      18'b000011011101010000: begin o_move = 4'd1; end
      18'b001100000100110101: begin o_move = 4'd1; end
      18'b001100011101010000: begin o_move = 4'd1; end
      18'b110000011101000100: begin o_move = 4'd2; end
      18'b110000011101010000: begin o_move = 4'd2; end
      18'b000000001101110101: begin o_move = 4'd3; end
      18'b001100000001110101: begin o_move = 4'd3; end
      18'b001100010000110101: begin o_move = 4'd3; end
      18'b110000011101000001: begin o_move = 4'd3; end
      18'b110100001101000001: begin o_move = 4'd3; end
      18'b110100001101000100: begin o_move = 4'd3; end
      18'b110111000001000100: begin o_move = 4'd5; end
      18'b110111000001010000: begin o_move = 4'd5; end
      18'b110111010000000001: begin o_move = 4'd5; end
      18'b110111010000000100: begin o_move = 4'd5; end
      18'b001101000000110101: begin o_move = 4'd6; end
      18'b110000011100000101: begin o_move = 4'd7; end
      18'b110001110101000000: begin o_move = 4'd7; end
      18'b110100001100000101: begin o_move = 4'd7; end
      18'b110100110101000000: begin o_move = 4'd7; end
      18'b110111000001000001: begin o_move = 4'd7; end
      18'b001101001100010001: begin o_move = 4'd8; end
      18'b001101001101010000: begin o_move = 4'd8; end
      18'b110000011100010001: begin o_move = 4'd8; end
      18'b110100001100010001: begin o_move = 4'd8; end
      18'b110111000100000001: begin o_move = 4'd8; end
      18'b110111000100010000: begin o_move = 4'd8; end
      18'b001101001100010100: begin o_move = 4'd9; end
      18'b110000011100010100: begin o_move = 4'd9; end
      18'b110100001100010100: begin o_move = 4'd9; end
      18'b110100001101010000: begin o_move = 4'd9; end
      18'b001101110101110100: begin o_move = 4'd1; end
      18'b000011011101011101: begin o_move = 4'd2; end
      18'b110000011101011101: begin o_move = 4'd2; end
      18'b110100001101011101: begin o_move = 4'd3; end
      18'b110111000100011101: begin o_move = 4'd4; end
      18'b110111000101001101: begin o_move = 4'd4; end
      18'b110111000101110001: begin o_move = 4'd4; end
      18'b110111010001110001: begin o_move = 4'd5; end
      18'b110111010100001101: begin o_move = 4'd6; end
      18'b110100110101001101: begin o_move = 4'd7; end
      18'b110111010111010000: begin o_move = 4'd9; end
      18'b001100011101110101: begin o_move = 4'd3; end
      18'b110000011101110101: begin o_move = 4'd3; end
      18'b110100001101110101: begin o_move = 4'd3; end
      18'b110111000001110101: begin o_move = 4'd4; end
      18'b110111011100000101: begin o_move = 4'd7; end
      18'b110111011101000001: begin o_move = 4'd7; end
      18'b110111011101000100: begin o_move = 4'd7; end
      18'b110111011100010001: begin o_move = 4'd8; end
      18'b110111011100010100: begin o_move = 4'd9; end
      18'b110111011101010000: begin o_move = 4'd9; end
      18'b110111001101000101: begin o_move = 4'd7; end
      18'b110111110101000001: begin o_move = 4'd7; end
      18'b110111001101010001: begin o_move = 4'd8; end
      18'b110111110101010000: begin o_move = 4'd8; end
      18'b110111001101010100: begin o_move = 4'd9; end
      18'b001111000101010111: begin o_move = 4'd1; end
      18'b001111010100010111: begin o_move = 4'd1; end
      18'b111100000101010111: begin o_move = 4'd3; end
      18'b111100010001010111: begin o_move = 4'd3; end
      18'b111100010100010111: begin o_move = 4'd3; end
      18'b111101000001010111: begin o_move = 4'd5; end
      18'b111101010000010111: begin o_move = 4'd5; end
      18'b000011110101000001: begin o_move = 4'd1; end
      18'b000011110101010000: begin o_move = 4'd1; end
      18'b000011110101000100: begin o_move = 4'd2; end
      18'b110000110101000100: begin o_move = 4'd2; end
      18'b110011000001000101: begin o_move = 4'd2; end
      18'b110011000001010001: begin o_move = 4'd2; end
      18'b110011000001010100: begin o_move = 4'd2; end
      18'b110011000100000101: begin o_move = 4'd2; end
      18'b110011000100010001: begin o_move = 4'd2; end
      18'b110011000100010100: begin o_move = 4'd2; end
      18'b110011000101000001: begin o_move = 4'd2; end
      18'b110011000101000100: begin o_move = 4'd2; end
      18'b110011000101010000: begin o_move = 4'd2; end
      18'b110011010000000101: begin o_move = 4'd2; end
      18'b110011010000010001: begin o_move = 4'd2; end
      18'b110011010000010100: begin o_move = 4'd2; end
      18'b110011010001000001: begin o_move = 4'd2; end
      18'b110011010001000100: begin o_move = 4'd2; end
      18'b110011010001010000: begin o_move = 4'd2; end
      18'b110011010100000001: begin o_move = 4'd2; end
      18'b110011010100000100: begin o_move = 4'd2; end
      18'b110011010100010000: begin o_move = 4'd2; end
      18'b110000110101000001: begin o_move = 4'd3; end
      18'b110000110101010000: begin o_move = 4'd3; end
      18'b111100000100000101: begin o_move = 4'd3; end
      18'b111100000100010100: begin o_move = 4'd3; end
      18'b111100000101000100: begin o_move = 4'd3; end
      18'b111100010000010001: begin o_move = 4'd3; end
      18'b111100010000010100: begin o_move = 4'd3; end
      18'b111100010001010000: begin o_move = 4'd3; end
      18'b111100010100000100: begin o_move = 4'd3; end
      18'b111100010100010000: begin o_move = 4'd3; end
      18'b111101010000010000: begin o_move = 4'd5; end
      18'b000011001101000101: begin o_move = 4'd7; end
      18'b111101000100000100: begin o_move = 4'd7; end
      18'b000011001101010001: begin o_move = 4'd8; end
      18'b001100001101010001: begin o_move = 4'd8; end
      18'b001100001101010100: begin o_move = 4'd9; end
      18'b111101000101110100: begin o_move = 4'd4; end
      18'b111101010100110100: begin o_move = 4'd6; end
      18'b111101010111000001: begin o_move = 4'd7; end
      18'b111101010111000100: begin o_move = 4'd7; end
      18'b001100110101110101: begin o_move = 4'd1; end
      18'b001111000101110101: begin o_move = 4'd1; end
      18'b001111010001110101: begin o_move = 4'd1; end
      18'b001111010100110101: begin o_move = 4'd1; end
      18'b110011010111010001: begin o_move = 4'd2; end
      18'b110011010111010100: begin o_move = 4'd2; end
      18'b111100000101110101: begin o_move = 4'd3; end
      18'b111100010100110101: begin o_move = 4'd3; end
      18'b111100010111000101: begin o_move = 4'd3; end
      18'b111100010111010001: begin o_move = 4'd3; end
      18'b111100010111010100: begin o_move = 4'd3; end
      18'b111101000100110101: begin o_move = 4'd4; end
      18'b111101011100010001: begin o_move = 4'd8; end
      18'b111101011101010000: begin o_move = 4'd8; end
      18'b111101011100010100: begin o_move = 4'd9; end
      18'b111101011101000100: begin o_move = 4'd9; end
      18'b110011011101000101: begin o_move = 4'd2; end
      18'b110011011101010001: begin o_move = 4'd2; end
      18'b110011011101010100: begin o_move = 4'd2; end
      18'b111100011101000101: begin o_move = 4'd3; end
      18'b111100011101010001: begin o_move = 4'd3; end
      18'b111100011101010100: begin o_move = 4'd3; end
      18'b111101110101000100: begin o_move = 4'd7; end
      18'b001111110101000101: begin o_move = 4'd1; end
      18'b001111110101010100: begin o_move = 4'd1; end
      18'b110011110101000101: begin o_move = 4'd2; end
      18'b110011110101010001: begin o_move = 4'd2; end
      18'b110011110101010100: begin o_move = 4'd2; end
      18'b111100110101000101: begin o_move = 4'd3; end
      18'b111100110101010100: begin o_move = 4'd3; end
      default: begin o_move = 4'd0; end	// Bad move
    endcase
endmodule
